magic
tech sky130A
magscale 1 2
timestamp 1685316190
<< obsli1 >>
rect 1104 2159 438840 437393
<< obsm1 >>
rect 934 76 439102 437424
<< metal2 >>
rect 16210 0 16266 800
rect 17038 0 17094 800
rect 17866 0 17922 800
rect 18694 0 18750 800
rect 19522 0 19578 800
rect 20350 0 20406 800
rect 21178 0 21234 800
rect 22006 0 22062 800
rect 22834 0 22890 800
rect 23662 0 23718 800
rect 24490 0 24546 800
rect 25318 0 25374 800
rect 26146 0 26202 800
rect 26974 0 27030 800
rect 27802 0 27858 800
rect 28630 0 28686 800
rect 29458 0 29514 800
rect 30286 0 30342 800
rect 31114 0 31170 800
rect 31942 0 31998 800
rect 32770 0 32826 800
rect 33598 0 33654 800
rect 34426 0 34482 800
rect 35254 0 35310 800
rect 36082 0 36138 800
rect 36910 0 36966 800
rect 37738 0 37794 800
rect 38566 0 38622 800
rect 39394 0 39450 800
rect 40222 0 40278 800
rect 41050 0 41106 800
rect 41878 0 41934 800
rect 42706 0 42762 800
rect 43534 0 43590 800
rect 44362 0 44418 800
rect 45190 0 45246 800
rect 46018 0 46074 800
rect 46846 0 46902 800
rect 47674 0 47730 800
rect 48502 0 48558 800
rect 49330 0 49386 800
rect 50158 0 50214 800
rect 50986 0 51042 800
rect 51814 0 51870 800
rect 52642 0 52698 800
rect 53470 0 53526 800
rect 54298 0 54354 800
rect 55126 0 55182 800
rect 55954 0 56010 800
rect 56782 0 56838 800
rect 57610 0 57666 800
rect 58438 0 58494 800
rect 59266 0 59322 800
rect 60094 0 60150 800
rect 60922 0 60978 800
rect 61750 0 61806 800
rect 62578 0 62634 800
rect 63406 0 63462 800
rect 64234 0 64290 800
rect 65062 0 65118 800
rect 65890 0 65946 800
rect 66718 0 66774 800
rect 67546 0 67602 800
rect 68374 0 68430 800
rect 69202 0 69258 800
rect 70030 0 70086 800
rect 70858 0 70914 800
rect 71686 0 71742 800
rect 72514 0 72570 800
rect 73342 0 73398 800
rect 74170 0 74226 800
rect 74998 0 75054 800
rect 75826 0 75882 800
rect 76654 0 76710 800
rect 77482 0 77538 800
rect 78310 0 78366 800
rect 79138 0 79194 800
rect 79966 0 80022 800
rect 80794 0 80850 800
rect 81622 0 81678 800
rect 82450 0 82506 800
rect 83278 0 83334 800
rect 84106 0 84162 800
rect 84934 0 84990 800
rect 85762 0 85818 800
rect 86590 0 86646 800
rect 87418 0 87474 800
rect 88246 0 88302 800
rect 89074 0 89130 800
rect 89902 0 89958 800
rect 90730 0 90786 800
rect 91558 0 91614 800
rect 92386 0 92442 800
rect 93214 0 93270 800
rect 94042 0 94098 800
rect 94870 0 94926 800
rect 95698 0 95754 800
rect 96526 0 96582 800
rect 97354 0 97410 800
rect 98182 0 98238 800
rect 99010 0 99066 800
rect 99838 0 99894 800
rect 100666 0 100722 800
rect 101494 0 101550 800
rect 102322 0 102378 800
rect 103150 0 103206 800
rect 103978 0 104034 800
rect 104806 0 104862 800
rect 105634 0 105690 800
rect 106462 0 106518 800
rect 107290 0 107346 800
rect 108118 0 108174 800
rect 108946 0 109002 800
rect 109774 0 109830 800
rect 110602 0 110658 800
rect 111430 0 111486 800
rect 112258 0 112314 800
rect 113086 0 113142 800
rect 113914 0 113970 800
rect 114742 0 114798 800
rect 115570 0 115626 800
rect 116398 0 116454 800
rect 117226 0 117282 800
rect 118054 0 118110 800
rect 118882 0 118938 800
rect 119710 0 119766 800
rect 120538 0 120594 800
rect 121366 0 121422 800
rect 122194 0 122250 800
rect 123022 0 123078 800
rect 123850 0 123906 800
rect 124678 0 124734 800
rect 125506 0 125562 800
rect 126334 0 126390 800
rect 127162 0 127218 800
rect 127990 0 128046 800
rect 128818 0 128874 800
rect 129646 0 129702 800
rect 130474 0 130530 800
rect 131302 0 131358 800
rect 132130 0 132186 800
rect 132958 0 133014 800
rect 133786 0 133842 800
rect 134614 0 134670 800
rect 135442 0 135498 800
rect 136270 0 136326 800
rect 137098 0 137154 800
rect 137926 0 137982 800
rect 138754 0 138810 800
rect 139582 0 139638 800
rect 140410 0 140466 800
rect 141238 0 141294 800
rect 142066 0 142122 800
rect 142894 0 142950 800
rect 143722 0 143778 800
rect 144550 0 144606 800
rect 145378 0 145434 800
rect 146206 0 146262 800
rect 147034 0 147090 800
rect 147862 0 147918 800
rect 148690 0 148746 800
rect 149518 0 149574 800
rect 150346 0 150402 800
rect 151174 0 151230 800
rect 152002 0 152058 800
rect 152830 0 152886 800
rect 153658 0 153714 800
rect 154486 0 154542 800
rect 155314 0 155370 800
rect 156142 0 156198 800
rect 156970 0 157026 800
rect 157798 0 157854 800
rect 158626 0 158682 800
rect 159454 0 159510 800
rect 160282 0 160338 800
rect 161110 0 161166 800
rect 161938 0 161994 800
rect 162766 0 162822 800
rect 163594 0 163650 800
rect 164422 0 164478 800
rect 165250 0 165306 800
rect 166078 0 166134 800
rect 166906 0 166962 800
rect 167734 0 167790 800
rect 168562 0 168618 800
rect 169390 0 169446 800
rect 170218 0 170274 800
rect 171046 0 171102 800
rect 171874 0 171930 800
rect 172702 0 172758 800
rect 173530 0 173586 800
rect 174358 0 174414 800
rect 175186 0 175242 800
rect 176014 0 176070 800
rect 176842 0 176898 800
rect 177670 0 177726 800
rect 178498 0 178554 800
rect 179326 0 179382 800
rect 180154 0 180210 800
rect 180982 0 181038 800
rect 181810 0 181866 800
rect 182638 0 182694 800
rect 183466 0 183522 800
rect 184294 0 184350 800
rect 185122 0 185178 800
rect 185950 0 186006 800
rect 186778 0 186834 800
rect 187606 0 187662 800
rect 188434 0 188490 800
rect 189262 0 189318 800
rect 190090 0 190146 800
rect 190918 0 190974 800
rect 191746 0 191802 800
rect 192574 0 192630 800
rect 193402 0 193458 800
rect 194230 0 194286 800
rect 195058 0 195114 800
rect 195886 0 195942 800
rect 196714 0 196770 800
rect 197542 0 197598 800
rect 198370 0 198426 800
rect 199198 0 199254 800
rect 200026 0 200082 800
rect 200854 0 200910 800
rect 201682 0 201738 800
rect 202510 0 202566 800
rect 203338 0 203394 800
rect 204166 0 204222 800
rect 204994 0 205050 800
rect 205822 0 205878 800
rect 206650 0 206706 800
rect 207478 0 207534 800
rect 208306 0 208362 800
rect 209134 0 209190 800
rect 209962 0 210018 800
rect 210790 0 210846 800
rect 211618 0 211674 800
rect 212446 0 212502 800
rect 213274 0 213330 800
rect 214102 0 214158 800
rect 214930 0 214986 800
rect 215758 0 215814 800
rect 216586 0 216642 800
rect 217414 0 217470 800
rect 218242 0 218298 800
rect 219070 0 219126 800
rect 219898 0 219954 800
rect 220726 0 220782 800
rect 221554 0 221610 800
rect 222382 0 222438 800
rect 223210 0 223266 800
rect 224038 0 224094 800
rect 224866 0 224922 800
rect 225694 0 225750 800
rect 226522 0 226578 800
rect 227350 0 227406 800
rect 228178 0 228234 800
rect 229006 0 229062 800
rect 229834 0 229890 800
rect 230662 0 230718 800
rect 231490 0 231546 800
rect 232318 0 232374 800
rect 233146 0 233202 800
rect 233974 0 234030 800
rect 234802 0 234858 800
rect 235630 0 235686 800
rect 236458 0 236514 800
rect 237286 0 237342 800
rect 238114 0 238170 800
rect 238942 0 238998 800
rect 239770 0 239826 800
rect 240598 0 240654 800
rect 241426 0 241482 800
rect 242254 0 242310 800
rect 243082 0 243138 800
rect 243910 0 243966 800
rect 244738 0 244794 800
rect 245566 0 245622 800
rect 246394 0 246450 800
rect 247222 0 247278 800
rect 248050 0 248106 800
rect 248878 0 248934 800
rect 249706 0 249762 800
rect 250534 0 250590 800
rect 251362 0 251418 800
rect 252190 0 252246 800
rect 253018 0 253074 800
rect 253846 0 253902 800
rect 254674 0 254730 800
rect 255502 0 255558 800
rect 256330 0 256386 800
rect 257158 0 257214 800
rect 257986 0 258042 800
rect 258814 0 258870 800
rect 259642 0 259698 800
rect 260470 0 260526 800
rect 261298 0 261354 800
rect 262126 0 262182 800
rect 262954 0 263010 800
rect 263782 0 263838 800
rect 264610 0 264666 800
rect 265438 0 265494 800
rect 266266 0 266322 800
rect 267094 0 267150 800
rect 267922 0 267978 800
rect 268750 0 268806 800
rect 269578 0 269634 800
rect 270406 0 270462 800
rect 271234 0 271290 800
rect 272062 0 272118 800
rect 272890 0 272946 800
rect 273718 0 273774 800
rect 274546 0 274602 800
rect 275374 0 275430 800
rect 276202 0 276258 800
rect 277030 0 277086 800
rect 277858 0 277914 800
rect 278686 0 278742 800
rect 279514 0 279570 800
rect 280342 0 280398 800
rect 281170 0 281226 800
rect 281998 0 282054 800
rect 282826 0 282882 800
rect 283654 0 283710 800
rect 284482 0 284538 800
rect 285310 0 285366 800
rect 286138 0 286194 800
rect 286966 0 287022 800
rect 287794 0 287850 800
rect 288622 0 288678 800
rect 289450 0 289506 800
rect 290278 0 290334 800
rect 291106 0 291162 800
rect 291934 0 291990 800
rect 292762 0 292818 800
rect 293590 0 293646 800
rect 294418 0 294474 800
rect 295246 0 295302 800
rect 296074 0 296130 800
rect 296902 0 296958 800
rect 297730 0 297786 800
rect 298558 0 298614 800
rect 299386 0 299442 800
rect 300214 0 300270 800
rect 301042 0 301098 800
rect 301870 0 301926 800
rect 302698 0 302754 800
rect 303526 0 303582 800
rect 304354 0 304410 800
rect 305182 0 305238 800
rect 306010 0 306066 800
rect 306838 0 306894 800
rect 307666 0 307722 800
rect 308494 0 308550 800
rect 309322 0 309378 800
rect 310150 0 310206 800
rect 310978 0 311034 800
rect 311806 0 311862 800
rect 312634 0 312690 800
rect 313462 0 313518 800
rect 314290 0 314346 800
rect 315118 0 315174 800
rect 315946 0 316002 800
rect 316774 0 316830 800
rect 317602 0 317658 800
rect 318430 0 318486 800
rect 319258 0 319314 800
rect 320086 0 320142 800
rect 320914 0 320970 800
rect 321742 0 321798 800
rect 322570 0 322626 800
rect 323398 0 323454 800
rect 324226 0 324282 800
rect 325054 0 325110 800
rect 325882 0 325938 800
rect 326710 0 326766 800
rect 327538 0 327594 800
rect 328366 0 328422 800
rect 329194 0 329250 800
rect 330022 0 330078 800
rect 330850 0 330906 800
rect 331678 0 331734 800
rect 332506 0 332562 800
rect 333334 0 333390 800
rect 334162 0 334218 800
rect 334990 0 335046 800
rect 335818 0 335874 800
rect 336646 0 336702 800
rect 337474 0 337530 800
rect 338302 0 338358 800
rect 339130 0 339186 800
rect 339958 0 340014 800
rect 340786 0 340842 800
rect 341614 0 341670 800
rect 342442 0 342498 800
rect 343270 0 343326 800
rect 344098 0 344154 800
rect 344926 0 344982 800
rect 345754 0 345810 800
rect 346582 0 346638 800
rect 347410 0 347466 800
rect 348238 0 348294 800
rect 349066 0 349122 800
rect 349894 0 349950 800
rect 350722 0 350778 800
rect 351550 0 351606 800
rect 352378 0 352434 800
rect 353206 0 353262 800
rect 354034 0 354090 800
rect 354862 0 354918 800
rect 355690 0 355746 800
rect 356518 0 356574 800
rect 357346 0 357402 800
rect 358174 0 358230 800
rect 359002 0 359058 800
rect 359830 0 359886 800
rect 360658 0 360714 800
rect 361486 0 361542 800
rect 362314 0 362370 800
rect 363142 0 363198 800
rect 363970 0 364026 800
rect 364798 0 364854 800
rect 365626 0 365682 800
rect 366454 0 366510 800
rect 367282 0 367338 800
rect 368110 0 368166 800
rect 368938 0 368994 800
rect 369766 0 369822 800
rect 370594 0 370650 800
rect 371422 0 371478 800
rect 372250 0 372306 800
rect 373078 0 373134 800
rect 373906 0 373962 800
rect 374734 0 374790 800
rect 375562 0 375618 800
rect 376390 0 376446 800
rect 377218 0 377274 800
rect 378046 0 378102 800
rect 378874 0 378930 800
rect 379702 0 379758 800
rect 380530 0 380586 800
rect 381358 0 381414 800
rect 382186 0 382242 800
rect 383014 0 383070 800
rect 383842 0 383898 800
rect 384670 0 384726 800
rect 385498 0 385554 800
rect 386326 0 386382 800
rect 387154 0 387210 800
rect 387982 0 388038 800
rect 388810 0 388866 800
rect 389638 0 389694 800
rect 390466 0 390522 800
rect 391294 0 391350 800
rect 392122 0 392178 800
rect 392950 0 393006 800
rect 393778 0 393834 800
rect 394606 0 394662 800
rect 395434 0 395490 800
rect 396262 0 396318 800
rect 397090 0 397146 800
rect 397918 0 397974 800
rect 398746 0 398802 800
rect 399574 0 399630 800
rect 400402 0 400458 800
rect 401230 0 401286 800
rect 402058 0 402114 800
rect 402886 0 402942 800
rect 403714 0 403770 800
rect 404542 0 404598 800
rect 405370 0 405426 800
rect 406198 0 406254 800
rect 407026 0 407082 800
rect 407854 0 407910 800
rect 408682 0 408738 800
rect 409510 0 409566 800
rect 410338 0 410394 800
rect 411166 0 411222 800
rect 411994 0 412050 800
rect 412822 0 412878 800
rect 413650 0 413706 800
rect 414478 0 414534 800
rect 415306 0 415362 800
rect 416134 0 416190 800
rect 416962 0 417018 800
rect 417790 0 417846 800
rect 418618 0 418674 800
rect 419446 0 419502 800
rect 420274 0 420330 800
rect 421102 0 421158 800
rect 421930 0 421986 800
rect 422758 0 422814 800
rect 423586 0 423642 800
<< obsm2 >>
rect 938 856 439098 437413
rect 938 70 16154 856
rect 16322 70 16982 856
rect 17150 70 17810 856
rect 17978 70 18638 856
rect 18806 70 19466 856
rect 19634 70 20294 856
rect 20462 70 21122 856
rect 21290 70 21950 856
rect 22118 70 22778 856
rect 22946 70 23606 856
rect 23774 70 24434 856
rect 24602 70 25262 856
rect 25430 70 26090 856
rect 26258 70 26918 856
rect 27086 70 27746 856
rect 27914 70 28574 856
rect 28742 70 29402 856
rect 29570 70 30230 856
rect 30398 70 31058 856
rect 31226 70 31886 856
rect 32054 70 32714 856
rect 32882 70 33542 856
rect 33710 70 34370 856
rect 34538 70 35198 856
rect 35366 70 36026 856
rect 36194 70 36854 856
rect 37022 70 37682 856
rect 37850 70 38510 856
rect 38678 70 39338 856
rect 39506 70 40166 856
rect 40334 70 40994 856
rect 41162 70 41822 856
rect 41990 70 42650 856
rect 42818 70 43478 856
rect 43646 70 44306 856
rect 44474 70 45134 856
rect 45302 70 45962 856
rect 46130 70 46790 856
rect 46958 70 47618 856
rect 47786 70 48446 856
rect 48614 70 49274 856
rect 49442 70 50102 856
rect 50270 70 50930 856
rect 51098 70 51758 856
rect 51926 70 52586 856
rect 52754 70 53414 856
rect 53582 70 54242 856
rect 54410 70 55070 856
rect 55238 70 55898 856
rect 56066 70 56726 856
rect 56894 70 57554 856
rect 57722 70 58382 856
rect 58550 70 59210 856
rect 59378 70 60038 856
rect 60206 70 60866 856
rect 61034 70 61694 856
rect 61862 70 62522 856
rect 62690 70 63350 856
rect 63518 70 64178 856
rect 64346 70 65006 856
rect 65174 70 65834 856
rect 66002 70 66662 856
rect 66830 70 67490 856
rect 67658 70 68318 856
rect 68486 70 69146 856
rect 69314 70 69974 856
rect 70142 70 70802 856
rect 70970 70 71630 856
rect 71798 70 72458 856
rect 72626 70 73286 856
rect 73454 70 74114 856
rect 74282 70 74942 856
rect 75110 70 75770 856
rect 75938 70 76598 856
rect 76766 70 77426 856
rect 77594 70 78254 856
rect 78422 70 79082 856
rect 79250 70 79910 856
rect 80078 70 80738 856
rect 80906 70 81566 856
rect 81734 70 82394 856
rect 82562 70 83222 856
rect 83390 70 84050 856
rect 84218 70 84878 856
rect 85046 70 85706 856
rect 85874 70 86534 856
rect 86702 70 87362 856
rect 87530 70 88190 856
rect 88358 70 89018 856
rect 89186 70 89846 856
rect 90014 70 90674 856
rect 90842 70 91502 856
rect 91670 70 92330 856
rect 92498 70 93158 856
rect 93326 70 93986 856
rect 94154 70 94814 856
rect 94982 70 95642 856
rect 95810 70 96470 856
rect 96638 70 97298 856
rect 97466 70 98126 856
rect 98294 70 98954 856
rect 99122 70 99782 856
rect 99950 70 100610 856
rect 100778 70 101438 856
rect 101606 70 102266 856
rect 102434 70 103094 856
rect 103262 70 103922 856
rect 104090 70 104750 856
rect 104918 70 105578 856
rect 105746 70 106406 856
rect 106574 70 107234 856
rect 107402 70 108062 856
rect 108230 70 108890 856
rect 109058 70 109718 856
rect 109886 70 110546 856
rect 110714 70 111374 856
rect 111542 70 112202 856
rect 112370 70 113030 856
rect 113198 70 113858 856
rect 114026 70 114686 856
rect 114854 70 115514 856
rect 115682 70 116342 856
rect 116510 70 117170 856
rect 117338 70 117998 856
rect 118166 70 118826 856
rect 118994 70 119654 856
rect 119822 70 120482 856
rect 120650 70 121310 856
rect 121478 70 122138 856
rect 122306 70 122966 856
rect 123134 70 123794 856
rect 123962 70 124622 856
rect 124790 70 125450 856
rect 125618 70 126278 856
rect 126446 70 127106 856
rect 127274 70 127934 856
rect 128102 70 128762 856
rect 128930 70 129590 856
rect 129758 70 130418 856
rect 130586 70 131246 856
rect 131414 70 132074 856
rect 132242 70 132902 856
rect 133070 70 133730 856
rect 133898 70 134558 856
rect 134726 70 135386 856
rect 135554 70 136214 856
rect 136382 70 137042 856
rect 137210 70 137870 856
rect 138038 70 138698 856
rect 138866 70 139526 856
rect 139694 70 140354 856
rect 140522 70 141182 856
rect 141350 70 142010 856
rect 142178 70 142838 856
rect 143006 70 143666 856
rect 143834 70 144494 856
rect 144662 70 145322 856
rect 145490 70 146150 856
rect 146318 70 146978 856
rect 147146 70 147806 856
rect 147974 70 148634 856
rect 148802 70 149462 856
rect 149630 70 150290 856
rect 150458 70 151118 856
rect 151286 70 151946 856
rect 152114 70 152774 856
rect 152942 70 153602 856
rect 153770 70 154430 856
rect 154598 70 155258 856
rect 155426 70 156086 856
rect 156254 70 156914 856
rect 157082 70 157742 856
rect 157910 70 158570 856
rect 158738 70 159398 856
rect 159566 70 160226 856
rect 160394 70 161054 856
rect 161222 70 161882 856
rect 162050 70 162710 856
rect 162878 70 163538 856
rect 163706 70 164366 856
rect 164534 70 165194 856
rect 165362 70 166022 856
rect 166190 70 166850 856
rect 167018 70 167678 856
rect 167846 70 168506 856
rect 168674 70 169334 856
rect 169502 70 170162 856
rect 170330 70 170990 856
rect 171158 70 171818 856
rect 171986 70 172646 856
rect 172814 70 173474 856
rect 173642 70 174302 856
rect 174470 70 175130 856
rect 175298 70 175958 856
rect 176126 70 176786 856
rect 176954 70 177614 856
rect 177782 70 178442 856
rect 178610 70 179270 856
rect 179438 70 180098 856
rect 180266 70 180926 856
rect 181094 70 181754 856
rect 181922 70 182582 856
rect 182750 70 183410 856
rect 183578 70 184238 856
rect 184406 70 185066 856
rect 185234 70 185894 856
rect 186062 70 186722 856
rect 186890 70 187550 856
rect 187718 70 188378 856
rect 188546 70 189206 856
rect 189374 70 190034 856
rect 190202 70 190862 856
rect 191030 70 191690 856
rect 191858 70 192518 856
rect 192686 70 193346 856
rect 193514 70 194174 856
rect 194342 70 195002 856
rect 195170 70 195830 856
rect 195998 70 196658 856
rect 196826 70 197486 856
rect 197654 70 198314 856
rect 198482 70 199142 856
rect 199310 70 199970 856
rect 200138 70 200798 856
rect 200966 70 201626 856
rect 201794 70 202454 856
rect 202622 70 203282 856
rect 203450 70 204110 856
rect 204278 70 204938 856
rect 205106 70 205766 856
rect 205934 70 206594 856
rect 206762 70 207422 856
rect 207590 70 208250 856
rect 208418 70 209078 856
rect 209246 70 209906 856
rect 210074 70 210734 856
rect 210902 70 211562 856
rect 211730 70 212390 856
rect 212558 70 213218 856
rect 213386 70 214046 856
rect 214214 70 214874 856
rect 215042 70 215702 856
rect 215870 70 216530 856
rect 216698 70 217358 856
rect 217526 70 218186 856
rect 218354 70 219014 856
rect 219182 70 219842 856
rect 220010 70 220670 856
rect 220838 70 221498 856
rect 221666 70 222326 856
rect 222494 70 223154 856
rect 223322 70 223982 856
rect 224150 70 224810 856
rect 224978 70 225638 856
rect 225806 70 226466 856
rect 226634 70 227294 856
rect 227462 70 228122 856
rect 228290 70 228950 856
rect 229118 70 229778 856
rect 229946 70 230606 856
rect 230774 70 231434 856
rect 231602 70 232262 856
rect 232430 70 233090 856
rect 233258 70 233918 856
rect 234086 70 234746 856
rect 234914 70 235574 856
rect 235742 70 236402 856
rect 236570 70 237230 856
rect 237398 70 238058 856
rect 238226 70 238886 856
rect 239054 70 239714 856
rect 239882 70 240542 856
rect 240710 70 241370 856
rect 241538 70 242198 856
rect 242366 70 243026 856
rect 243194 70 243854 856
rect 244022 70 244682 856
rect 244850 70 245510 856
rect 245678 70 246338 856
rect 246506 70 247166 856
rect 247334 70 247994 856
rect 248162 70 248822 856
rect 248990 70 249650 856
rect 249818 70 250478 856
rect 250646 70 251306 856
rect 251474 70 252134 856
rect 252302 70 252962 856
rect 253130 70 253790 856
rect 253958 70 254618 856
rect 254786 70 255446 856
rect 255614 70 256274 856
rect 256442 70 257102 856
rect 257270 70 257930 856
rect 258098 70 258758 856
rect 258926 70 259586 856
rect 259754 70 260414 856
rect 260582 70 261242 856
rect 261410 70 262070 856
rect 262238 70 262898 856
rect 263066 70 263726 856
rect 263894 70 264554 856
rect 264722 70 265382 856
rect 265550 70 266210 856
rect 266378 70 267038 856
rect 267206 70 267866 856
rect 268034 70 268694 856
rect 268862 70 269522 856
rect 269690 70 270350 856
rect 270518 70 271178 856
rect 271346 70 272006 856
rect 272174 70 272834 856
rect 273002 70 273662 856
rect 273830 70 274490 856
rect 274658 70 275318 856
rect 275486 70 276146 856
rect 276314 70 276974 856
rect 277142 70 277802 856
rect 277970 70 278630 856
rect 278798 70 279458 856
rect 279626 70 280286 856
rect 280454 70 281114 856
rect 281282 70 281942 856
rect 282110 70 282770 856
rect 282938 70 283598 856
rect 283766 70 284426 856
rect 284594 70 285254 856
rect 285422 70 286082 856
rect 286250 70 286910 856
rect 287078 70 287738 856
rect 287906 70 288566 856
rect 288734 70 289394 856
rect 289562 70 290222 856
rect 290390 70 291050 856
rect 291218 70 291878 856
rect 292046 70 292706 856
rect 292874 70 293534 856
rect 293702 70 294362 856
rect 294530 70 295190 856
rect 295358 70 296018 856
rect 296186 70 296846 856
rect 297014 70 297674 856
rect 297842 70 298502 856
rect 298670 70 299330 856
rect 299498 70 300158 856
rect 300326 70 300986 856
rect 301154 70 301814 856
rect 301982 70 302642 856
rect 302810 70 303470 856
rect 303638 70 304298 856
rect 304466 70 305126 856
rect 305294 70 305954 856
rect 306122 70 306782 856
rect 306950 70 307610 856
rect 307778 70 308438 856
rect 308606 70 309266 856
rect 309434 70 310094 856
rect 310262 70 310922 856
rect 311090 70 311750 856
rect 311918 70 312578 856
rect 312746 70 313406 856
rect 313574 70 314234 856
rect 314402 70 315062 856
rect 315230 70 315890 856
rect 316058 70 316718 856
rect 316886 70 317546 856
rect 317714 70 318374 856
rect 318542 70 319202 856
rect 319370 70 320030 856
rect 320198 70 320858 856
rect 321026 70 321686 856
rect 321854 70 322514 856
rect 322682 70 323342 856
rect 323510 70 324170 856
rect 324338 70 324998 856
rect 325166 70 325826 856
rect 325994 70 326654 856
rect 326822 70 327482 856
rect 327650 70 328310 856
rect 328478 70 329138 856
rect 329306 70 329966 856
rect 330134 70 330794 856
rect 330962 70 331622 856
rect 331790 70 332450 856
rect 332618 70 333278 856
rect 333446 70 334106 856
rect 334274 70 334934 856
rect 335102 70 335762 856
rect 335930 70 336590 856
rect 336758 70 337418 856
rect 337586 70 338246 856
rect 338414 70 339074 856
rect 339242 70 339902 856
rect 340070 70 340730 856
rect 340898 70 341558 856
rect 341726 70 342386 856
rect 342554 70 343214 856
rect 343382 70 344042 856
rect 344210 70 344870 856
rect 345038 70 345698 856
rect 345866 70 346526 856
rect 346694 70 347354 856
rect 347522 70 348182 856
rect 348350 70 349010 856
rect 349178 70 349838 856
rect 350006 70 350666 856
rect 350834 70 351494 856
rect 351662 70 352322 856
rect 352490 70 353150 856
rect 353318 70 353978 856
rect 354146 70 354806 856
rect 354974 70 355634 856
rect 355802 70 356462 856
rect 356630 70 357290 856
rect 357458 70 358118 856
rect 358286 70 358946 856
rect 359114 70 359774 856
rect 359942 70 360602 856
rect 360770 70 361430 856
rect 361598 70 362258 856
rect 362426 70 363086 856
rect 363254 70 363914 856
rect 364082 70 364742 856
rect 364910 70 365570 856
rect 365738 70 366398 856
rect 366566 70 367226 856
rect 367394 70 368054 856
rect 368222 70 368882 856
rect 369050 70 369710 856
rect 369878 70 370538 856
rect 370706 70 371366 856
rect 371534 70 372194 856
rect 372362 70 373022 856
rect 373190 70 373850 856
rect 374018 70 374678 856
rect 374846 70 375506 856
rect 375674 70 376334 856
rect 376502 70 377162 856
rect 377330 70 377990 856
rect 378158 70 378818 856
rect 378986 70 379646 856
rect 379814 70 380474 856
rect 380642 70 381302 856
rect 381470 70 382130 856
rect 382298 70 382958 856
rect 383126 70 383786 856
rect 383954 70 384614 856
rect 384782 70 385442 856
rect 385610 70 386270 856
rect 386438 70 387098 856
rect 387266 70 387926 856
rect 388094 70 388754 856
rect 388922 70 389582 856
rect 389750 70 390410 856
rect 390578 70 391238 856
rect 391406 70 392066 856
rect 392234 70 392894 856
rect 393062 70 393722 856
rect 393890 70 394550 856
rect 394718 70 395378 856
rect 395546 70 396206 856
rect 396374 70 397034 856
rect 397202 70 397862 856
rect 398030 70 398690 856
rect 398858 70 399518 856
rect 399686 70 400346 856
rect 400514 70 401174 856
rect 401342 70 402002 856
rect 402170 70 402830 856
rect 402998 70 403658 856
rect 403826 70 404486 856
rect 404654 70 405314 856
rect 405482 70 406142 856
rect 406310 70 406970 856
rect 407138 70 407798 856
rect 407966 70 408626 856
rect 408794 70 409454 856
rect 409622 70 410282 856
rect 410450 70 411110 856
rect 411278 70 411938 856
rect 412106 70 412766 856
rect 412934 70 413594 856
rect 413762 70 414422 856
rect 414590 70 415250 856
rect 415418 70 416078 856
rect 416246 70 416906 856
rect 417074 70 417734 856
rect 417902 70 418562 856
rect 418730 70 419390 856
rect 419558 70 420218 856
rect 420386 70 421046 856
rect 421214 70 421874 856
rect 422042 70 422702 856
rect 422870 70 423530 856
rect 423698 70 439098 856
<< metal3 >>
rect 0 433168 800 433288
rect 439200 433168 440000 433288
rect 0 425552 800 425672
rect 439200 425552 440000 425672
rect 0 417936 800 418056
rect 439200 417936 440000 418056
rect 0 410320 800 410440
rect 439200 410320 440000 410440
rect 0 402704 800 402824
rect 439200 402704 440000 402824
rect 0 395088 800 395208
rect 439200 395088 440000 395208
rect 0 387472 800 387592
rect 439200 387472 440000 387592
rect 0 379856 800 379976
rect 439200 379856 440000 379976
rect 0 372240 800 372360
rect 439200 372240 440000 372360
rect 0 364624 800 364744
rect 439200 364624 440000 364744
rect 0 357008 800 357128
rect 439200 357008 440000 357128
rect 0 349392 800 349512
rect 439200 349392 440000 349512
rect 0 341776 800 341896
rect 439200 341776 440000 341896
rect 0 334160 800 334280
rect 439200 334160 440000 334280
rect 0 326544 800 326664
rect 439200 326544 440000 326664
rect 0 318928 800 319048
rect 439200 318928 440000 319048
rect 0 311312 800 311432
rect 439200 311312 440000 311432
rect 0 303696 800 303816
rect 439200 303696 440000 303816
rect 0 296080 800 296200
rect 439200 296080 440000 296200
rect 0 288464 800 288584
rect 439200 288464 440000 288584
rect 0 280848 800 280968
rect 439200 280848 440000 280968
rect 0 273232 800 273352
rect 439200 273232 440000 273352
rect 0 265616 800 265736
rect 439200 265616 440000 265736
rect 0 258000 800 258120
rect 439200 258000 440000 258120
rect 0 250384 800 250504
rect 439200 250384 440000 250504
rect 0 242768 800 242888
rect 439200 242768 440000 242888
rect 0 235152 800 235272
rect 439200 235152 440000 235272
rect 0 227536 800 227656
rect 439200 227536 440000 227656
rect 0 219920 800 220040
rect 439200 219920 440000 220040
rect 0 212304 800 212424
rect 439200 212304 440000 212424
rect 0 204688 800 204808
rect 439200 204688 440000 204808
rect 0 197072 800 197192
rect 439200 197072 440000 197192
rect 0 189456 800 189576
rect 439200 189456 440000 189576
rect 0 181840 800 181960
rect 439200 181840 440000 181960
rect 0 174224 800 174344
rect 439200 174224 440000 174344
rect 0 166608 800 166728
rect 439200 166608 440000 166728
rect 0 158992 800 159112
rect 439200 158992 440000 159112
rect 0 151376 800 151496
rect 439200 151376 440000 151496
rect 0 143760 800 143880
rect 439200 143760 440000 143880
rect 0 136144 800 136264
rect 439200 136144 440000 136264
rect 0 128528 800 128648
rect 439200 128528 440000 128648
rect 0 120912 800 121032
rect 439200 120912 440000 121032
rect 0 113296 800 113416
rect 439200 113296 440000 113416
rect 0 105680 800 105800
rect 439200 105680 440000 105800
rect 0 98064 800 98184
rect 439200 98064 440000 98184
rect 0 90448 800 90568
rect 439200 90448 440000 90568
rect 0 82832 800 82952
rect 439200 82832 440000 82952
rect 0 75216 800 75336
rect 439200 75216 440000 75336
rect 0 67600 800 67720
rect 439200 67600 440000 67720
rect 0 59984 800 60104
rect 439200 59984 440000 60104
rect 0 52368 800 52488
rect 439200 52368 440000 52488
rect 0 44752 800 44872
rect 439200 44752 440000 44872
rect 0 37136 800 37256
rect 439200 37136 440000 37256
rect 0 29520 800 29640
rect 439200 29520 440000 29640
rect 0 21904 800 22024
rect 439200 21904 440000 22024
rect 0 14288 800 14408
rect 439200 14288 440000 14408
rect 0 6672 800 6792
rect 439200 6672 440000 6792
<< obsm3 >>
rect 800 433368 439200 437409
rect 880 433088 439120 433368
rect 800 425752 439200 433088
rect 880 425472 439120 425752
rect 800 418136 439200 425472
rect 880 417856 439120 418136
rect 800 410520 439200 417856
rect 880 410240 439120 410520
rect 800 402904 439200 410240
rect 880 402624 439120 402904
rect 800 395288 439200 402624
rect 880 395008 439120 395288
rect 800 387672 439200 395008
rect 880 387392 439120 387672
rect 800 380056 439200 387392
rect 880 379776 439120 380056
rect 800 372440 439200 379776
rect 880 372160 439120 372440
rect 800 364824 439200 372160
rect 880 364544 439120 364824
rect 800 357208 439200 364544
rect 880 356928 439120 357208
rect 800 349592 439200 356928
rect 880 349312 439120 349592
rect 800 341976 439200 349312
rect 880 341696 439120 341976
rect 800 334360 439200 341696
rect 880 334080 439120 334360
rect 800 326744 439200 334080
rect 880 326464 439120 326744
rect 800 319128 439200 326464
rect 880 318848 439120 319128
rect 800 311512 439200 318848
rect 880 311232 439120 311512
rect 800 303896 439200 311232
rect 880 303616 439120 303896
rect 800 296280 439200 303616
rect 880 296000 439120 296280
rect 800 288664 439200 296000
rect 880 288384 439120 288664
rect 800 281048 439200 288384
rect 880 280768 439120 281048
rect 800 273432 439200 280768
rect 880 273152 439120 273432
rect 800 265816 439200 273152
rect 880 265536 439120 265816
rect 800 258200 439200 265536
rect 880 257920 439120 258200
rect 800 250584 439200 257920
rect 880 250304 439120 250584
rect 800 242968 439200 250304
rect 880 242688 439120 242968
rect 800 235352 439200 242688
rect 880 235072 439120 235352
rect 800 227736 439200 235072
rect 880 227456 439120 227736
rect 800 220120 439200 227456
rect 880 219840 439120 220120
rect 800 212504 439200 219840
rect 880 212224 439120 212504
rect 800 204888 439200 212224
rect 880 204608 439120 204888
rect 800 197272 439200 204608
rect 880 196992 439120 197272
rect 800 189656 439200 196992
rect 880 189376 439120 189656
rect 800 182040 439200 189376
rect 880 181760 439120 182040
rect 800 174424 439200 181760
rect 880 174144 439120 174424
rect 800 166808 439200 174144
rect 880 166528 439120 166808
rect 800 159192 439200 166528
rect 880 158912 439120 159192
rect 800 151576 439200 158912
rect 880 151296 439120 151576
rect 800 143960 439200 151296
rect 880 143680 439120 143960
rect 800 136344 439200 143680
rect 880 136064 439120 136344
rect 800 128728 439200 136064
rect 880 128448 439120 128728
rect 800 121112 439200 128448
rect 880 120832 439120 121112
rect 800 113496 439200 120832
rect 880 113216 439120 113496
rect 800 105880 439200 113216
rect 880 105600 439120 105880
rect 800 98264 439200 105600
rect 880 97984 439120 98264
rect 800 90648 439200 97984
rect 880 90368 439120 90648
rect 800 83032 439200 90368
rect 880 82752 439120 83032
rect 800 75416 439200 82752
rect 880 75136 439120 75416
rect 800 67800 439200 75136
rect 880 67520 439120 67800
rect 800 60184 439200 67520
rect 880 59904 439120 60184
rect 800 52568 439200 59904
rect 880 52288 439120 52568
rect 800 44952 439200 52288
rect 880 44672 439120 44952
rect 800 37336 439200 44672
rect 880 37056 439120 37336
rect 800 29720 439200 37056
rect 880 29440 439120 29720
rect 800 22104 439200 29440
rect 880 21824 439120 22104
rect 800 14488 439200 21824
rect 880 14208 439120 14488
rect 800 6872 439200 14208
rect 880 6592 439120 6872
rect 800 307 439200 6592
<< metal4 >>
rect 4208 2128 4528 437424
rect 19568 2128 19888 437424
rect 34928 2128 35248 437424
rect 50288 2128 50608 437424
rect 65648 2128 65968 437424
rect 81008 2128 81328 437424
rect 96368 2128 96688 437424
rect 111728 2128 112048 437424
rect 127088 2128 127408 437424
rect 142448 2128 142768 437424
rect 157808 2128 158128 437424
rect 173168 2128 173488 437424
rect 188528 2128 188848 437424
rect 203888 2128 204208 437424
rect 219248 2128 219568 437424
rect 234608 2128 234928 437424
rect 249968 2128 250288 437424
rect 265328 2128 265648 437424
rect 280688 2128 281008 437424
rect 296048 2128 296368 437424
rect 311408 2128 311728 437424
rect 326768 2128 327088 437424
rect 342128 2128 342448 437424
rect 357488 2128 357808 437424
rect 372848 2128 373168 437424
rect 388208 2128 388528 437424
rect 403568 2128 403888 437424
rect 418928 2128 419248 437424
rect 434288 2128 434608 437424
<< obsm4 >>
rect 127939 2048 142368 417485
rect 142848 2048 157728 417485
rect 158208 2048 173088 417485
rect 173568 2048 188448 417485
rect 188928 2048 203808 417485
rect 204288 2048 219168 417485
rect 219648 2048 234528 417485
rect 235008 2048 249888 417485
rect 250368 2048 265248 417485
rect 265728 2048 280608 417485
rect 281088 2048 295968 417485
rect 296448 2048 311328 417485
rect 311808 2048 326688 417485
rect 327168 2048 342048 417485
rect 342528 2048 357408 417485
rect 357888 2048 372768 417485
rect 373248 2048 388128 417485
rect 388608 2048 403488 417485
rect 403968 2048 418848 417485
rect 419328 2048 434208 417485
rect 434688 2048 436573 417485
rect 127939 443 436573 2048
<< labels >>
rlabel metal3 s 439200 6672 440000 6792 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 439200 235152 440000 235272 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 439200 258000 440000 258120 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 439200 280848 440000 280968 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 439200 303696 440000 303816 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 439200 326544 440000 326664 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 439200 349392 440000 349512 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 439200 372240 440000 372360 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 439200 395088 440000 395208 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 439200 417936 440000 418056 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 433168 800 433288 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 439200 29520 440000 29640 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 410320 800 410440 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 387472 800 387592 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 364624 800 364744 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 341776 800 341896 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 318928 800 319048 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 296080 800 296200 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 273232 800 273352 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 250384 800 250504 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 227536 800 227656 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 204688 800 204808 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 439200 52368 440000 52488 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 181840 800 181960 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 158992 800 159112 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 136144 800 136264 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 113296 800 113416 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 439200 75216 440000 75336 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 439200 98064 440000 98184 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 439200 120912 440000 121032 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 439200 143760 440000 143880 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 439200 166608 440000 166728 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 439200 189456 440000 189576 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 439200 212304 440000 212424 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 439200 21904 440000 22024 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 439200 250384 440000 250504 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 439200 273232 440000 273352 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 439200 296080 440000 296200 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 439200 318928 440000 319048 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 439200 341776 440000 341896 6 io_oeb[14]
port 44 nsew signal output
rlabel metal3 s 439200 364624 440000 364744 6 io_oeb[15]
port 45 nsew signal output
rlabel metal3 s 439200 387472 440000 387592 6 io_oeb[16]
port 46 nsew signal output
rlabel metal3 s 439200 410320 440000 410440 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 439200 433168 440000 433288 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 417936 800 418056 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 439200 44752 440000 44872 6 io_oeb[1]
port 50 nsew signal output
rlabel metal3 s 0 395088 800 395208 6 io_oeb[20]
port 51 nsew signal output
rlabel metal3 s 0 372240 800 372360 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 0 349392 800 349512 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 0 326544 800 326664 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 303696 800 303816 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 280848 800 280968 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 258000 800 258120 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 235152 800 235272 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 212304 800 212424 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 189456 800 189576 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 439200 67600 440000 67720 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 166608 800 166728 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 143760 800 143880 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 120912 800 121032 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 98064 800 98184 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 75216 800 75336 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 439200 90448 440000 90568 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 439200 113296 440000 113416 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 439200 136144 440000 136264 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 439200 158992 440000 159112 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 439200 181840 440000 181960 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 439200 204688 440000 204808 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 439200 227536 440000 227656 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 439200 14288 440000 14408 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 439200 242768 440000 242888 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 439200 265616 440000 265736 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 439200 288464 440000 288584 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 439200 311312 440000 311432 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 439200 334160 440000 334280 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 439200 357008 440000 357128 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 439200 379856 440000 379976 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 439200 402704 440000 402824 6 io_out[17]
port 85 nsew signal output
rlabel metal3 s 439200 425552 440000 425672 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 0 425552 800 425672 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 439200 37136 440000 37256 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 0 402704 800 402824 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 0 379856 800 379976 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 0 357008 800 357128 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 0 334160 800 334280 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 311312 800 311432 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 288464 800 288584 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 265616 800 265736 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 242768 800 242888 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 219920 800 220040 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 197072 800 197192 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 439200 59984 440000 60104 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 174224 800 174344 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 151376 800 151496 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 128528 800 128648 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 105680 800 105800 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 82832 800 82952 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 59984 800 60104 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 439200 82832 440000 82952 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 439200 105680 440000 105800 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 439200 128528 440000 128648 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 439200 151376 440000 151496 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 439200 174224 440000 174344 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 439200 197072 440000 197192 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 439200 219920 440000 220040 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 421930 0 421986 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 422758 0 422814 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 423586 0 423642 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 352378 0 352434 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 354862 0 354918 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 357346 0 357402 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 359830 0 359886 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 362314 0 362370 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 364798 0 364854 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 367282 0 367338 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 369766 0 369822 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 372250 0 372306 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 374734 0 374790 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 377218 0 377274 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 379702 0 379758 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 382186 0 382242 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 384670 0 384726 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 387154 0 387210 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 389638 0 389694 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 392122 0 392178 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 394606 0 394662 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 397090 0 397146 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 399574 0 399630 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 402058 0 402114 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 404542 0 404598 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 407026 0 407082 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 409510 0 409566 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 411994 0 412050 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 414478 0 414534 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 416962 0 417018 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 419446 0 419502 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 166078 0 166134 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 176014 0 176070 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 178498 0 178554 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 185950 0 186006 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 188434 0 188490 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 190918 0 190974 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 193402 0 193458 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 195886 0 195942 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 198370 0 198426 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 200854 0 200910 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 203338 0 203394 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 205822 0 205878 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 208306 0 208362 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 210790 0 210846 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 213274 0 213330 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 220726 0 220782 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 223210 0 223266 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 228178 0 228234 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 230662 0 230718 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 233146 0 233202 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 238114 0 238170 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 240598 0 240654 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 243082 0 243138 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 248050 0 248106 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 250534 0 250590 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 253018 0 253074 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 255502 0 255558 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 257986 0 258042 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 260470 0 260526 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 262954 0 263010 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 265438 0 265494 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 267922 0 267978 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 270406 0 270462 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 272890 0 272946 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 275374 0 275430 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 277858 0 277914 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 280342 0 280398 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 282826 0 282882 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 285310 0 285366 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 287794 0 287850 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 290278 0 290334 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 292762 0 292818 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 295246 0 295302 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 297730 0 297786 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 300214 0 300270 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 302698 0 302754 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 305182 0 305238 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 307666 0 307722 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 310150 0 310206 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 312634 0 312690 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 315118 0 315174 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 317602 0 317658 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 320086 0 320142 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 322570 0 322626 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 325054 0 325110 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 327538 0 327594 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 330022 0 330078 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 332506 0 332562 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 334990 0 335046 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 337474 0 337530 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 339958 0 340014 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 342442 0 342498 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 344926 0 344982 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 347410 0 347466 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 349894 0 349950 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 353206 0 353262 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 355690 0 355746 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 358174 0 358230 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 360658 0 360714 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 363142 0 363198 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 365626 0 365682 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 368110 0 368166 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 370594 0 370650 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 373078 0 373134 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 375562 0 375618 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 129646 0 129702 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 378046 0 378102 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 380530 0 380586 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 383014 0 383070 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 385498 0 385554 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 387982 0 388038 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 390466 0 390522 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 392950 0 393006 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 395434 0 395490 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 397918 0 397974 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 400402 0 400458 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 402886 0 402942 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 405370 0 405426 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 407854 0 407910 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 410338 0 410394 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 412822 0 412878 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 415306 0 415362 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 417790 0 417846 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 420274 0 420330 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 137098 0 137154 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 142066 0 142122 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 144550 0 144606 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 154486 0 154542 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 159454 0 159510 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 164422 0 164478 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 169390 0 169446 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 171874 0 171930 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 179326 0 179382 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 181810 0 181866 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 184294 0 184350 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 186778 0 186834 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 189262 0 189318 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 191746 0 191802 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 194230 0 194286 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 196714 0 196770 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 199198 0 199254 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 201682 0 201738 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 206650 0 206706 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 209134 0 209190 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 211618 0 211674 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 214102 0 214158 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 216586 0 216642 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 219070 0 219126 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 221554 0 221610 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 224038 0 224094 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 226522 0 226578 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 114742 0 114798 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 229006 0 229062 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 231490 0 231546 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 233974 0 234030 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 236458 0 236514 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 238942 0 238998 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 241426 0 241482 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 243910 0 243966 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 246394 0 246450 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 248878 0 248934 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 251362 0 251418 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 253846 0 253902 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 256330 0 256386 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 258814 0 258870 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 261298 0 261354 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 263782 0 263838 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 266266 0 266322 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 268750 0 268806 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 271234 0 271290 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 273718 0 273774 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 276202 0 276258 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 278686 0 278742 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 281170 0 281226 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 283654 0 283710 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 286138 0 286194 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 288622 0 288678 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 291106 0 291162 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 293590 0 293646 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 296074 0 296130 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 298558 0 298614 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 301042 0 301098 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 122194 0 122250 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 303526 0 303582 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 306010 0 306066 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 308494 0 308550 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 310978 0 311034 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 313462 0 313518 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 315946 0 316002 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 318430 0 318486 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 320914 0 320970 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 323398 0 323454 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 325882 0 325938 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 328366 0 328422 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 330850 0 330906 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 333334 0 333390 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 335818 0 335874 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 338302 0 338358 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 340786 0 340842 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 343270 0 343326 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 345754 0 345810 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 348238 0 348294 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 350722 0 350778 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 354034 0 354090 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 356518 0 356574 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 359002 0 359058 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 361486 0 361542 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 363970 0 364026 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 366454 0 366510 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 368938 0 368994 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 371422 0 371478 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 373906 0 373962 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 376390 0 376446 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 378874 0 378930 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 381358 0 381414 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 383842 0 383898 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 386326 0 386382 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 388810 0 388866 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 391294 0 391350 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 393778 0 393834 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 396262 0 396318 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 398746 0 398802 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 401230 0 401286 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 403714 0 403770 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 406198 0 406254 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 408682 0 408738 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 411166 0 411222 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 413650 0 413706 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 416134 0 416190 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 418618 0 418674 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 421102 0 421158 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 165250 0 165306 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 172702 0 172758 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 180154 0 180210 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 185122 0 185178 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 187606 0 187662 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 190090 0 190146 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 200026 0 200082 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 202510 0 202566 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 204994 0 205050 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 207478 0 207534 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 209962 0 210018 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 212446 0 212502 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 214930 0 214986 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 217414 0 217470 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 219898 0 219954 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 222382 0 222438 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 224866 0 224922 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 227350 0 227406 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 229834 0 229890 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 232318 0 232374 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 234802 0 234858 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 237286 0 237342 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 239770 0 239826 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 242254 0 242310 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 244738 0 244794 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 247222 0 247278 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 249706 0 249762 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 252190 0 252246 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 254674 0 254730 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 257158 0 257214 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 259642 0 259698 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 262126 0 262182 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 264610 0 264666 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 267094 0 267150 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 269578 0 269634 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 272062 0 272118 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 274546 0 274602 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 277030 0 277086 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 279514 0 279570 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 281998 0 282054 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 284482 0 284538 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 286966 0 287022 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 289450 0 289506 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 291934 0 291990 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 294418 0 294474 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 296902 0 296958 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 299386 0 299442 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 301870 0 301926 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 304354 0 304410 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 306838 0 306894 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 309322 0 309378 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 311806 0 311862 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 314290 0 314346 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 316774 0 316830 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 319258 0 319314 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 321742 0 321798 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 324226 0 324282 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 326710 0 326766 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 329194 0 329250 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 331678 0 331734 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 334162 0 334218 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 336646 0 336702 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 339130 0 339186 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 341614 0 341670 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 344098 0 344154 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 346582 0 346638 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 349066 0 349122 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 351550 0 351606 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 16210 0 16266 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 78310 0 78366 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 103150 0 103206 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 440000 440000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 171013068
string GDS_FILE /ux1/users/asinghan/18224-tapeout-s23-caravel/openlane/user_proj/runs/23_05_28_17_40/results/signoff/user_proj.magic.gds
string GDS_START 1936512
<< end >>

